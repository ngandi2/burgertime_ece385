// /*
//  * ECE385-HelperTools/PNG-To-Txt
//  * Author: Rishi Thakkar
//  *
//  */

// module spriteRAM
// (
// 	input [4:0] data_In,
// 	input [18:0] write_address, read_address,
// 	input we, Clk,
// 	output logic [4:0] data_Out
// );

// // mem has width of 3 bits and a total of 42240 addresses
// // ['0x000000', '0xFF0000', '0xFFFFFF', '0x6D6D6D', '0xFFFF00', '0x00FF00', '0xFFB600', '0x6DB600']
// logic [2:0] mem [0:42239];

// initial
// begin
// 	 $readmemh("sprite_bytes/sprites.txt", mem);
// end


// always_ff @ (posedge Clk) begin
// 	if (we)
// 		mem[write_address] <= data_In;
// 	data_Out<= mem[read_address];
// end

// endmodule
